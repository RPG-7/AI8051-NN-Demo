module sdram_controller_top #(

);



endmodule

